`include "../databook/gates.v"
`include "../circuit.v"

module ALU(y, a, b, cin);


module MicroWaveRange(clk1, clk2, r, p);
    input clk1, clk2, r, p;
